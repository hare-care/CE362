module multiply(
    input clk, rstn,
    input [31:0],
    output []
);

endmodule